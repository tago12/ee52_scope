-- sopc_scope_sys.vhd

-- Generated using ACDS version 13.1 162 at 2014.04.25.21:41:18

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sopc_scope_sys is
	port (
		clk_clk                             : in    std_logic                     := '0';             --        clk.clk
		bridge_out_addr_out                 : out   std_logic_vector(18 downto 0);                    -- bridge_out.addr_out
		bridge_out_rom_tcm_chipselect_n_out : out   std_logic_vector(0 downto 0);                     --           .rom_tcm_chipselect_n_out
		bridge_out_ram_tcm_read_out         : out   std_logic_vector(0 downto 0);                     --           .ram_tcm_read_out
		bridge_out_ram_tcm_write_n_out      : out   std_logic_vector(0 downto 0);                     --           .ram_tcm_write_n_out
		bridge_out_data_outen               : inout std_logic_vector(7 downto 0)  := (others => '0'); --           .data_outen
		bridge_out_rom_tcm_read_out         : out   std_logic_vector(0 downto 0);                     --           .rom_tcm_read_out
		bridge_out_ram_tcm_chipselect_n_out : out   std_logic_vector(0 downto 0)                      --           .ram_tcm_chipselect_n_out
	);
end entity sopc_scope_sys;

architecture rtl of sopc_scope_sys is
	component sopc_scope_sys_nios is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(20 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(20 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component sopc_scope_sys_nios;

	component sopc_scope_sys_temp_ram is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(7 downto 0);                     -- readdata
			writedata  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component sopc_scope_sys_temp_ram;

	component sopc_scope_sys_jtag is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component sopc_scope_sys_jtag;

	component sopc_scope_sys_ram is
		generic (
			TCM_ADDRESS_W                  : integer := 30;
			TCM_DATA_W                     : integer := 32;
			TCM_BYTEENABLE_W               : integer := 4;
			TCM_READ_WAIT                  : integer := 1;
			TCM_WRITE_WAIT                 : integer := 0;
			TCM_SETUP_WAIT                 : integer := 0;
			TCM_DATA_HOLD                  : integer := 0;
			TCM_TURNAROUND_TIME            : integer := 2;
			TCM_TIMING_UNITS               : integer := 1;
			TCM_READLATENCY                : integer := 2;
			TCM_SYMBOLS_PER_WORD           : integer := 4;
			USE_READDATA                   : integer := 1;
			USE_WRITEDATA                  : integer := 1;
			USE_READ                       : integer := 1;
			USE_WRITE                      : integer := 1;
			USE_BYTEENABLE                 : integer := 1;
			USE_CHIPSELECT                 : integer := 0;
			USE_LOCK                       : integer := 0;
			USE_ADDRESS                    : integer := 1;
			USE_WAITREQUEST                : integer := 0;
			USE_WRITEBYTEENABLE            : integer := 0;
			USE_OUTPUTENABLE               : integer := 0;
			USE_RESETREQUEST               : integer := 0;
			USE_IRQ                        : integer := 0;
			USE_RESET_OUTPUT               : integer := 0;
			ACTIVE_LOW_READ                : integer := 0;
			ACTIVE_LOW_LOCK                : integer := 0;
			ACTIVE_LOW_WRITE               : integer := 0;
			ACTIVE_LOW_CHIPSELECT          : integer := 0;
			ACTIVE_LOW_BYTEENABLE          : integer := 0;
			ACTIVE_LOW_OUTPUTENABLE        : integer := 0;
			ACTIVE_LOW_WRITEBYTEENABLE     : integer := 0;
			ACTIVE_LOW_WAITREQUEST         : integer := 0;
			ACTIVE_LOW_BEGINTRANSFER       : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			reset_reset          : in  std_logic                     := 'X';             -- reset
			uas_address          : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			uas_burstcount       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			uas_read             : in  std_logic                     := 'X';             -- read
			uas_write            : in  std_logic                     := 'X';             -- write
			uas_waitrequest      : out std_logic;                                        -- waitrequest
			uas_readdatavalid    : out std_logic;                                        -- readdatavalid
			uas_byteenable       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- byteenable
			uas_readdata         : out std_logic_vector(7 downto 0);                     -- readdata
			uas_writedata        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			uas_lock             : in  std_logic                     := 'X';             -- lock
			uas_debugaccess      : in  std_logic                     := 'X';             -- debugaccess
			tcm_write_n_out      : out std_logic;                                        -- write_n_out
			tcm_read_out         : out std_logic;                                        -- read_out
			tcm_chipselect_n_out : out std_logic;                                        -- chipselect_n_out
			tcm_request          : out std_logic;                                        -- request
			tcm_grant            : in  std_logic                     := 'X';             -- grant
			tcm_address_out      : out std_logic_vector(16 downto 0);                    -- address_out
			tcm_data_out         : out std_logic_vector(7 downto 0);                     -- data_out
			tcm_data_outen       : out std_logic;                                        -- data_outen
			tcm_data_in          : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- data_in
		);
	end component sopc_scope_sys_ram;

	component sopc_scope_sys_pin_sharer is
		port (
			clk_clk                  : in  std_logic                     := 'X';             -- clk
			reset_reset              : in  std_logic                     := 'X';             -- reset
			request                  : out std_logic;                                        -- request
			grant                    : in  std_logic                     := 'X';             -- grant
			rom_tcm_read_out         : out std_logic_vector(0 downto 0);                     -- rom_tcm_read_out_out
			rom_tcm_chipselect_n_out : out std_logic_vector(0 downto 0);                     -- rom_tcm_chipselect_n_out_out
			ram_tcm_write_n_out      : out std_logic_vector(0 downto 0);                     -- ram_tcm_write_n_out_out
			ram_tcm_read_out         : out std_logic_vector(0 downto 0);                     -- ram_tcm_read_out_out
			ram_tcm_chipselect_n_out : out std_logic_vector(0 downto 0);                     -- ram_tcm_chipselect_n_out_out
			addr_out                 : out std_logic_vector(18 downto 0);                    -- addr_out_out
			data_outen               : out std_logic_vector(7 downto 0);                     -- data_outen_out
			data_outen_in            : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- data_outen_in
			data_outen_outen         : out std_logic;                                        -- data_outen_outen
			tcs0_request             : in  std_logic                     := 'X';             -- request
			tcs0_grant               : out std_logic;                                        -- grant
			tcs0_address_out         : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address_out
			tcs0_write_n_out         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- write_n_out
			tcs0_read_out            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- read_out
			tcs0_data_out            : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- data_out
			tcs0_data_in             : out std_logic_vector(7 downto 0);                     -- data_in
			tcs0_data_outen          : in  std_logic                     := 'X';             -- data_outen
			tcs0_chipselect_n_out    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- chipselect_n_out
			tcs1_request             : in  std_logic                     := 'X';             -- request
			tcs1_grant               : out std_logic;                                        -- grant
			tcs1_address_out         : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address_out
			tcs1_read_out            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- read_out
			tcs1_data_out            : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- data_out
			tcs1_data_in             : out std_logic_vector(7 downto 0);                     -- data_in
			tcs1_data_outen          : in  std_logic                     := 'X';             -- data_outen
			tcs1_chipselect_n_out    : in  std_logic_vector(0 downto 0)  := (others => 'X')  -- chipselect_n_out
		);
	end component sopc_scope_sys_pin_sharer;

	component sopc_scope_sys_bridge is
		port (
			clk                          : in    std_logic                     := 'X';             -- clk
			reset                        : in    std_logic                     := 'X';             -- reset
			request                      : in    std_logic                     := 'X';             -- request
			grant                        : out   std_logic;                                        -- grant
			tcs_addr_out                 : in    std_logic_vector(18 downto 0) := (others => 'X'); -- addr_out_out
			tcs_rom_tcm_chipselect_n_out : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- rom_tcm_chipselect_n_out_out
			tcs_ram_tcm_read_out         : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- ram_tcm_read_out_out
			tcs_ram_tcm_write_n_out      : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- ram_tcm_write_n_out_out
			tcs_data_outen               : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- data_outen_out
			tcs_data_outen_outen         : in    std_logic                     := 'X';             -- data_outen_outen
			tcs_data_outen_in            : out   std_logic_vector(7 downto 0);                     -- data_outen_in
			tcs_rom_tcm_read_out         : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- rom_tcm_read_out_out
			tcs_ram_tcm_chipselect_n_out : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- ram_tcm_chipselect_n_out_out
			addr_out                     : out   std_logic_vector(18 downto 0);                    -- addr_out
			rom_tcm_chipselect_n_out     : out   std_logic_vector(0 downto 0);                     -- rom_tcm_chipselect_n_out
			ram_tcm_read_out             : out   std_logic_vector(0 downto 0);                     -- ram_tcm_read_out
			ram_tcm_write_n_out          : out   std_logic_vector(0 downto 0);                     -- ram_tcm_write_n_out
			data_outen                   : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- data_outen
			rom_tcm_read_out             : out   std_logic_vector(0 downto 0);                     -- rom_tcm_read_out
			ram_tcm_chipselect_n_out     : out   std_logic_vector(0 downto 0)                      -- ram_tcm_chipselect_n_out
		);
	end component sopc_scope_sys_bridge;

	component sopc_scope_sys_rom is
		generic (
			TCM_ADDRESS_W                  : integer := 30;
			TCM_DATA_W                     : integer := 32;
			TCM_BYTEENABLE_W               : integer := 4;
			TCM_READ_WAIT                  : integer := 1;
			TCM_WRITE_WAIT                 : integer := 0;
			TCM_SETUP_WAIT                 : integer := 0;
			TCM_DATA_HOLD                  : integer := 0;
			TCM_TURNAROUND_TIME            : integer := 2;
			TCM_TIMING_UNITS               : integer := 1;
			TCM_READLATENCY                : integer := 2;
			TCM_SYMBOLS_PER_WORD           : integer := 4;
			USE_READDATA                   : integer := 1;
			USE_WRITEDATA                  : integer := 1;
			USE_READ                       : integer := 1;
			USE_WRITE                      : integer := 1;
			USE_BYTEENABLE                 : integer := 1;
			USE_CHIPSELECT                 : integer := 0;
			USE_LOCK                       : integer := 0;
			USE_ADDRESS                    : integer := 1;
			USE_WAITREQUEST                : integer := 0;
			USE_WRITEBYTEENABLE            : integer := 0;
			USE_OUTPUTENABLE               : integer := 0;
			USE_RESETREQUEST               : integer := 0;
			USE_IRQ                        : integer := 0;
			USE_RESET_OUTPUT               : integer := 0;
			ACTIVE_LOW_READ                : integer := 0;
			ACTIVE_LOW_LOCK                : integer := 0;
			ACTIVE_LOW_WRITE               : integer := 0;
			ACTIVE_LOW_CHIPSELECT          : integer := 0;
			ACTIVE_LOW_BYTEENABLE          : integer := 0;
			ACTIVE_LOW_OUTPUTENABLE        : integer := 0;
			ACTIVE_LOW_WRITEBYTEENABLE     : integer := 0;
			ACTIVE_LOW_WAITREQUEST         : integer := 0;
			ACTIVE_LOW_BEGINTRANSFER       : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			reset_reset          : in  std_logic                     := 'X';             -- reset
			uas_address          : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			uas_burstcount       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			uas_read             : in  std_logic                     := 'X';             -- read
			uas_write            : in  std_logic                     := 'X';             -- write
			uas_waitrequest      : out std_logic;                                        -- waitrequest
			uas_readdatavalid    : out std_logic;                                        -- readdatavalid
			uas_byteenable       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- byteenable
			uas_readdata         : out std_logic_vector(7 downto 0);                     -- readdata
			uas_writedata        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			uas_lock             : in  std_logic                     := 'X';             -- lock
			uas_debugaccess      : in  std_logic                     := 'X';             -- debugaccess
			tcm_read_out         : out std_logic;                                        -- read_out
			tcm_chipselect_n_out : out std_logic;                                        -- chipselect_n_out
			tcm_request          : out std_logic;                                        -- request
			tcm_grant            : in  std_logic                     := 'X';             -- grant
			tcm_address_out      : out std_logic_vector(18 downto 0);                    -- address_out
			tcm_data_out         : out std_logic_vector(7 downto 0);                     -- data_out
			tcm_data_outen       : out std_logic;                                        -- data_outen
			tcm_data_in          : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- data_in
		);
	end component sopc_scope_sys_rom;

	component sopc_scope_sys_mm_interconnect_0 is
		port (
			clk_0_clk_clk                            : in  std_logic                     := 'X';             -- clk
			nios_reset_n_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios_data_master_address                 : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			nios_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			nios_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios_data_master_read                    : in  std_logic                     := 'X';             -- read
			nios_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			nios_data_master_readdatavalid           : out std_logic;                                        -- readdatavalid
			nios_data_master_write                   : in  std_logic                     := 'X';             -- write
			nios_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			nios_instruction_master_address          : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			nios_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			nios_instruction_master_read             : in  std_logic                     := 'X';             -- read
			nios_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			nios_instruction_master_readdatavalid    : out std_logic;                                        -- readdatavalid
			jtag_avalon_jtag_slave_address           : out std_logic_vector(0 downto 0);                     -- address
			jtag_avalon_jtag_slave_write             : out std_logic;                                        -- write
			jtag_avalon_jtag_slave_read              : out std_logic;                                        -- read
			jtag_avalon_jtag_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_avalon_jtag_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_avalon_jtag_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			jtag_avalon_jtag_slave_chipselect        : out std_logic;                                        -- chipselect
			nios_jtag_debug_module_address           : out std_logic_vector(8 downto 0);                     -- address
			nios_jtag_debug_module_write             : out std_logic;                                        -- write
			nios_jtag_debug_module_read              : out std_logic;                                        -- read
			nios_jtag_debug_module_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios_jtag_debug_module_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios_jtag_debug_module_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios_jtag_debug_module_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios_jtag_debug_module_debugaccess       : out std_logic;                                        -- debugaccess
			ram_uas_address                          : out std_logic_vector(16 downto 0);                    -- address
			ram_uas_write                            : out std_logic;                                        -- write
			ram_uas_read                             : out std_logic;                                        -- read
			ram_uas_readdata                         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			ram_uas_writedata                        : out std_logic_vector(7 downto 0);                     -- writedata
			ram_uas_burstcount                       : out std_logic_vector(0 downto 0);                     -- burstcount
			ram_uas_byteenable                       : out std_logic_vector(0 downto 0);                     -- byteenable
			ram_uas_readdatavalid                    : in  std_logic                     := 'X';             -- readdatavalid
			ram_uas_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			ram_uas_lock                             : out std_logic;                                        -- lock
			ram_uas_debugaccess                      : out std_logic;                                        -- debugaccess
			rom_uas_address                          : out std_logic_vector(18 downto 0);                    -- address
			rom_uas_write                            : out std_logic;                                        -- write
			rom_uas_read                             : out std_logic;                                        -- read
			rom_uas_readdata                         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			rom_uas_writedata                        : out std_logic_vector(7 downto 0);                     -- writedata
			rom_uas_burstcount                       : out std_logic_vector(0 downto 0);                     -- burstcount
			rom_uas_byteenable                       : out std_logic_vector(0 downto 0);                     -- byteenable
			rom_uas_readdatavalid                    : in  std_logic                     := 'X';             -- readdatavalid
			rom_uas_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			rom_uas_lock                             : out std_logic;                                        -- lock
			rom_uas_debugaccess                      : out std_logic;                                        -- debugaccess
			temp_ram_s1_address                      : out std_logic_vector(15 downto 0);                    -- address
			temp_ram_s1_write                        : out std_logic;                                        -- write
			temp_ram_s1_readdata                     : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			temp_ram_s1_writedata                    : out std_logic_vector(7 downto 0);                     -- writedata
			temp_ram_s1_chipselect                   : out std_logic;                                        -- chipselect
			temp_ram_s1_clken                        : out std_logic                                         -- clken
		);
	end component sopc_scope_sys_mm_interconnect_0;

	component sopc_scope_sys_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component sopc_scope_sys_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal nios_jtag_debug_module_reset_reset                       : std_logic;                     -- nios:jtag_debug_module_resetrequest -> [rst_controller:reset_in0, rst_controller:reset_in1]
	signal ram_tcm_chipselect_n_out                                 : std_logic;                     -- ram:tcm_chipselect_n_out -> pin_sharer:tcs0_chipselect_n_out
	signal ram_tcm_grant                                            : std_logic;                     -- pin_sharer:tcs0_grant -> ram:tcm_grant
	signal ram_tcm_data_outen                                       : std_logic;                     -- ram:tcm_data_outen -> pin_sharer:tcs0_data_outen
	signal ram_tcm_request                                          : std_logic;                     -- ram:tcm_request -> pin_sharer:tcs0_request
	signal ram_tcm_data_out                                         : std_logic_vector(7 downto 0);  -- ram:tcm_data_out -> pin_sharer:tcs0_data_out
	signal ram_tcm_write_n_out                                      : std_logic;                     -- ram:tcm_write_n_out -> pin_sharer:tcs0_write_n_out
	signal ram_tcm_address_out                                      : std_logic_vector(16 downto 0); -- ram:tcm_address_out -> pin_sharer:tcs0_address_out
	signal ram_tcm_data_in                                          : std_logic_vector(7 downto 0);  -- pin_sharer:tcs0_data_in -> ram:tcm_data_in
	signal ram_tcm_read_out                                         : std_logic;                     -- ram:tcm_read_out -> pin_sharer:tcs0_read_out
	signal pin_sharer_tcm_rom_tcm_read_out_out                      : std_logic_vector(0 downto 0);  -- pin_sharer:rom_tcm_read_out -> bridge:tcs_rom_tcm_read_out
	signal pin_sharer_tcm_data_outen_outen                          : std_logic;                     -- pin_sharer:data_outen_outen -> bridge:tcs_data_outen_outen
	signal pin_sharer_tcm_addr_out_out                              : std_logic_vector(18 downto 0); -- pin_sharer:addr_out -> bridge:tcs_addr_out
	signal pin_sharer_tcm_data_outen_out                            : std_logic_vector(7 downto 0);  -- pin_sharer:data_outen -> bridge:tcs_data_outen
	signal pin_sharer_tcm_ram_tcm_chipselect_n_out_out              : std_logic_vector(0 downto 0);  -- pin_sharer:ram_tcm_chipselect_n_out -> bridge:tcs_ram_tcm_chipselect_n_out
	signal pin_sharer_tcm_grant                                     : std_logic;                     -- bridge:grant -> pin_sharer:grant
	signal pin_sharer_tcm_rom_tcm_chipselect_n_out_out              : std_logic_vector(0 downto 0);  -- pin_sharer:rom_tcm_chipselect_n_out -> bridge:tcs_rom_tcm_chipselect_n_out
	signal pin_sharer_tcm_request                                   : std_logic;                     -- pin_sharer:request -> bridge:request
	signal pin_sharer_tcm_data_outen_in                             : std_logic_vector(7 downto 0);  -- bridge:tcs_data_outen_in -> pin_sharer:data_outen_in
	signal pin_sharer_tcm_ram_tcm_write_n_out_out                   : std_logic_vector(0 downto 0);  -- pin_sharer:ram_tcm_write_n_out -> bridge:tcs_ram_tcm_write_n_out
	signal pin_sharer_tcm_ram_tcm_read_out_out                      : std_logic_vector(0 downto 0);  -- pin_sharer:ram_tcm_read_out -> bridge:tcs_ram_tcm_read_out
	signal rom_tcm_chipselect_n_out                                 : std_logic;                     -- rom:tcm_chipselect_n_out -> pin_sharer:tcs1_chipselect_n_out
	signal rom_tcm_grant                                            : std_logic;                     -- pin_sharer:tcs1_grant -> rom:tcm_grant
	signal rom_tcm_data_outen                                       : std_logic;                     -- rom:tcm_data_outen -> pin_sharer:tcs1_data_outen
	signal rom_tcm_request                                          : std_logic;                     -- rom:tcm_request -> pin_sharer:tcs1_request
	signal rom_tcm_data_out                                         : std_logic_vector(7 downto 0);  -- rom:tcm_data_out -> pin_sharer:tcs1_data_out
	signal rom_tcm_address_out                                      : std_logic_vector(18 downto 0); -- rom:tcm_address_out -> pin_sharer:tcs1_address_out
	signal rom_tcm_data_in                                          : std_logic_vector(7 downto 0);  -- pin_sharer:tcs1_data_in -> rom:tcm_data_in
	signal rom_tcm_read_out                                         : std_logic;                     -- rom:tcm_read_out -> pin_sharer:tcs1_read_out
	signal nios_data_master_waitrequest                             : std_logic;                     -- mm_interconnect_0:nios_data_master_waitrequest -> nios:d_waitrequest
	signal nios_data_master_writedata                               : std_logic_vector(31 downto 0); -- nios:d_writedata -> mm_interconnect_0:nios_data_master_writedata
	signal nios_data_master_address                                 : std_logic_vector(20 downto 0); -- nios:d_address -> mm_interconnect_0:nios_data_master_address
	signal nios_data_master_write                                   : std_logic;                     -- nios:d_write -> mm_interconnect_0:nios_data_master_write
	signal nios_data_master_read                                    : std_logic;                     -- nios:d_read -> mm_interconnect_0:nios_data_master_read
	signal nios_data_master_readdata                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_data_master_readdata -> nios:d_readdata
	signal nios_data_master_debugaccess                             : std_logic;                     -- nios:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios_data_master_debugaccess
	signal nios_data_master_readdatavalid                           : std_logic;                     -- mm_interconnect_0:nios_data_master_readdatavalid -> nios:d_readdatavalid
	signal nios_data_master_byteenable                              : std_logic_vector(3 downto 0);  -- nios:d_byteenable -> mm_interconnect_0:nios_data_master_byteenable
	signal mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	signal mm_interconnect_0_jtag_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	signal mm_interconnect_0_jtag_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	signal mm_interconnect_0_jtag_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_avalon_jtag_slave_write -> mm_interconnect_0_jtag_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_avalon_jtag_slave_read -> mm_interconnect_0_jtag_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	signal mm_interconnect_0_ram_uas_waitrequest                    : std_logic;                     -- ram:uas_waitrequest -> mm_interconnect_0:ram_uas_waitrequest
	signal mm_interconnect_0_ram_uas_burstcount                     : std_logic_vector(0 downto 0);  -- mm_interconnect_0:ram_uas_burstcount -> ram:uas_burstcount
	signal mm_interconnect_0_ram_uas_writedata                      : std_logic_vector(7 downto 0);  -- mm_interconnect_0:ram_uas_writedata -> ram:uas_writedata
	signal mm_interconnect_0_ram_uas_address                        : std_logic_vector(16 downto 0); -- mm_interconnect_0:ram_uas_address -> ram:uas_address
	signal mm_interconnect_0_ram_uas_lock                           : std_logic;                     -- mm_interconnect_0:ram_uas_lock -> ram:uas_lock
	signal mm_interconnect_0_ram_uas_write                          : std_logic;                     -- mm_interconnect_0:ram_uas_write -> ram:uas_write
	signal mm_interconnect_0_ram_uas_read                           : std_logic;                     -- mm_interconnect_0:ram_uas_read -> ram:uas_read
	signal mm_interconnect_0_ram_uas_readdata                       : std_logic_vector(7 downto 0);  -- ram:uas_readdata -> mm_interconnect_0:ram_uas_readdata
	signal mm_interconnect_0_ram_uas_debugaccess                    : std_logic;                     -- mm_interconnect_0:ram_uas_debugaccess -> ram:uas_debugaccess
	signal mm_interconnect_0_ram_uas_readdatavalid                  : std_logic;                     -- ram:uas_readdatavalid -> mm_interconnect_0:ram_uas_readdatavalid
	signal mm_interconnect_0_ram_uas_byteenable                     : std_logic_vector(0 downto 0);  -- mm_interconnect_0:ram_uas_byteenable -> ram:uas_byteenable
	signal mm_interconnect_0_rom_uas_waitrequest                    : std_logic;                     -- rom:uas_waitrequest -> mm_interconnect_0:rom_uas_waitrequest
	signal mm_interconnect_0_rom_uas_burstcount                     : std_logic_vector(0 downto 0);  -- mm_interconnect_0:rom_uas_burstcount -> rom:uas_burstcount
	signal mm_interconnect_0_rom_uas_writedata                      : std_logic_vector(7 downto 0);  -- mm_interconnect_0:rom_uas_writedata -> rom:uas_writedata
	signal mm_interconnect_0_rom_uas_address                        : std_logic_vector(18 downto 0); -- mm_interconnect_0:rom_uas_address -> rom:uas_address
	signal mm_interconnect_0_rom_uas_lock                           : std_logic;                     -- mm_interconnect_0:rom_uas_lock -> rom:uas_lock
	signal mm_interconnect_0_rom_uas_write                          : std_logic;                     -- mm_interconnect_0:rom_uas_write -> rom:uas_write
	signal mm_interconnect_0_rom_uas_read                           : std_logic;                     -- mm_interconnect_0:rom_uas_read -> rom:uas_read
	signal mm_interconnect_0_rom_uas_readdata                       : std_logic_vector(7 downto 0);  -- rom:uas_readdata -> mm_interconnect_0:rom_uas_readdata
	signal mm_interconnect_0_rom_uas_debugaccess                    : std_logic;                     -- mm_interconnect_0:rom_uas_debugaccess -> rom:uas_debugaccess
	signal mm_interconnect_0_rom_uas_readdatavalid                  : std_logic;                     -- rom:uas_readdatavalid -> mm_interconnect_0:rom_uas_readdatavalid
	signal mm_interconnect_0_rom_uas_byteenable                     : std_logic_vector(0 downto 0);  -- mm_interconnect_0:rom_uas_byteenable -> rom:uas_byteenable
	signal mm_interconnect_0_temp_ram_s1_writedata                  : std_logic_vector(7 downto 0);  -- mm_interconnect_0:temp_ram_s1_writedata -> temp_ram:writedata
	signal mm_interconnect_0_temp_ram_s1_address                    : std_logic_vector(15 downto 0); -- mm_interconnect_0:temp_ram_s1_address -> temp_ram:address
	signal mm_interconnect_0_temp_ram_s1_chipselect                 : std_logic;                     -- mm_interconnect_0:temp_ram_s1_chipselect -> temp_ram:chipselect
	signal mm_interconnect_0_temp_ram_s1_clken                      : std_logic;                     -- mm_interconnect_0:temp_ram_s1_clken -> temp_ram:clken
	signal mm_interconnect_0_temp_ram_s1_write                      : std_logic;                     -- mm_interconnect_0:temp_ram_s1_write -> temp_ram:write
	signal mm_interconnect_0_temp_ram_s1_readdata                   : std_logic_vector(7 downto 0);  -- temp_ram:readdata -> mm_interconnect_0:temp_ram_s1_readdata
	signal nios_instruction_master_waitrequest                      : std_logic;                     -- mm_interconnect_0:nios_instruction_master_waitrequest -> nios:i_waitrequest
	signal nios_instruction_master_address                          : std_logic_vector(20 downto 0); -- nios:i_address -> mm_interconnect_0:nios_instruction_master_address
	signal nios_instruction_master_read                             : std_logic;                     -- nios:i_read -> mm_interconnect_0:nios_instruction_master_read
	signal nios_instruction_master_readdata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_instruction_master_readdata -> nios:i_readdata
	signal nios_instruction_master_readdatavalid                    : std_logic;                     -- mm_interconnect_0:nios_instruction_master_readdatavalid -> nios:i_readdatavalid
	signal mm_interconnect_0_nios_jtag_debug_module_waitrequest     : std_logic;                     -- nios:jtag_debug_module_waitrequest -> mm_interconnect_0:nios_jtag_debug_module_waitrequest
	signal mm_interconnect_0_nios_jtag_debug_module_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_jtag_debug_module_writedata -> nios:jtag_debug_module_writedata
	signal mm_interconnect_0_nios_jtag_debug_module_address         : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios_jtag_debug_module_address -> nios:jtag_debug_module_address
	signal mm_interconnect_0_nios_jtag_debug_module_write           : std_logic;                     -- mm_interconnect_0:nios_jtag_debug_module_write -> nios:jtag_debug_module_write
	signal mm_interconnect_0_nios_jtag_debug_module_read            : std_logic;                     -- mm_interconnect_0:nios_jtag_debug_module_read -> nios:jtag_debug_module_read
	signal mm_interconnect_0_nios_jtag_debug_module_readdata        : std_logic_vector(31 downto 0); -- nios:jtag_debug_module_readdata -> mm_interconnect_0:nios_jtag_debug_module_readdata
	signal mm_interconnect_0_nios_jtag_debug_module_debugaccess     : std_logic;                     -- mm_interconnect_0:nios_jtag_debug_module_debugaccess -> nios:jtag_debug_module_debugaccess
	signal mm_interconnect_0_nios_jtag_debug_module_byteenable      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios_jtag_debug_module_byteenable -> nios:jtag_debug_module_byteenable
	signal irq_mapper_receiver0_irq                                 : std_logic;                     -- jtag:av_irq -> irq_mapper:receiver0_irq
	signal nios_d_irq_irq                                           : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios:d_irq
	signal rst_controller_reset_out_reset                           : std_logic;                     -- rst_controller:reset_out -> [bridge:reset, irq_mapper:reset, mm_interconnect_0:nios_reset_n_reset_bridge_in_reset_reset, pin_sharer:reset_reset, ram:reset_reset, rom:reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset, temp_ram:reset]
	signal rst_controller_reset_out_reset_req                       : std_logic;                     -- rst_controller:reset_req -> [nios:reset_req, rst_translator:reset_req_in, temp_ram:reset_req]
	signal mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_avalon_jtag_slave_write:inv -> jtag:av_write_n
	signal mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_avalon_jtag_slave_read:inv -> jtag:av_read_n
	signal rst_controller_reset_out_reset_ports_inv                 : std_logic;                     -- rst_controller_reset_out_reset:inv -> [jtag:rst_n, nios:reset_n]

begin

	nios : component sopc_scope_sys_nios
		port map (
			clk                                   => clk_clk,                                              --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,             --                   reset_n.reset_n
			reset_req                             => rst_controller_reset_out_reset_req,                   --                          .reset_req
			d_address                             => nios_data_master_address,                             --               data_master.address
			d_byteenable                          => nios_data_master_byteenable,                          --                          .byteenable
			d_read                                => nios_data_master_read,                                --                          .read
			d_readdata                            => nios_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => nios_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => nios_data_master_write,                               --                          .write
			d_writedata                           => nios_data_master_writedata,                           --                          .writedata
			d_readdatavalid                       => nios_data_master_readdatavalid,                       --                          .readdatavalid
			jtag_debug_module_debugaccess_to_roms => nios_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => nios_instruction_master_address,                      --        instruction_master.address
			i_read                                => nios_instruction_master_read,                         --                          .read
			i_readdata                            => nios_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => nios_instruction_master_waitrequest,                  --                          .waitrequest
			i_readdatavalid                       => nios_instruction_master_readdatavalid,                --                          .readdatavalid
			d_irq                                 => nios_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => nios_jtag_debug_module_reset_reset,                   --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_0_nios_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_0_nios_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_0_nios_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_0_nios_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_0_nios_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_0_nios_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_0_nios_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_0_nios_jtag_debug_module_writedata,   --                          .writedata
			no_ci_readra                          => open                                                  -- custom_instruction_master.readra
		);

	temp_ram : component sopc_scope_sys_temp_ram
		port map (
			clk        => clk_clk,                                  --   clk1.clk
			address    => mm_interconnect_0_temp_ram_s1_address,    --     s1.address
			clken      => mm_interconnect_0_temp_ram_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_temp_ram_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_temp_ram_s1_write,      --       .write
			readdata   => mm_interconnect_0_temp_ram_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_temp_ram_s1_writedata,  --       .writedata
			reset      => rst_controller_reset_out_reset,           -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req        --       .reset_req
		);

	jtag : component sopc_scope_sys_jtag
		port map (
			clk            => clk_clk,                                                  --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                 --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                  --               irq.irq
		);

	ram : component sopc_scope_sys_ram
		generic map (
			TCM_ADDRESS_W                  => 17,
			TCM_DATA_W                     => 8,
			TCM_BYTEENABLE_W               => 1,
			TCM_READ_WAIT                  => 3,
			TCM_WRITE_WAIT                 => 3,
			TCM_SETUP_WAIT                 => 0,
			TCM_DATA_HOLD                  => 1,
			TCM_TURNAROUND_TIME            => 2,
			TCM_TIMING_UNITS               => 1,
			TCM_READLATENCY                => 2,
			TCM_SYMBOLS_PER_WORD           => 1,
			USE_READDATA                   => 1,
			USE_WRITEDATA                  => 1,
			USE_READ                       => 1,
			USE_WRITE                      => 1,
			USE_BYTEENABLE                 => 0,
			USE_CHIPSELECT                 => 1,
			USE_LOCK                       => 0,
			USE_ADDRESS                    => 1,
			USE_WAITREQUEST                => 0,
			USE_WRITEBYTEENABLE            => 0,
			USE_OUTPUTENABLE               => 0,
			USE_RESETREQUEST               => 0,
			USE_IRQ                        => 0,
			USE_RESET_OUTPUT               => 0,
			ACTIVE_LOW_READ                => 0,
			ACTIVE_LOW_LOCK                => 0,
			ACTIVE_LOW_WRITE               => 1,
			ACTIVE_LOW_CHIPSELECT          => 1,
			ACTIVE_LOW_BYTEENABLE          => 0,
			ACTIVE_LOW_OUTPUTENABLE        => 0,
			ACTIVE_LOW_WRITEBYTEENABLE     => 0,
			ACTIVE_LOW_WAITREQUEST         => 0,
			ACTIVE_LOW_BEGINTRANSFER       => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0
		)
		port map (
			clk_clk              => clk_clk,                                 --   clk.clk
			reset_reset          => rst_controller_reset_out_reset,          -- reset.reset
			uas_address          => mm_interconnect_0_ram_uas_address,       --   uas.address
			uas_burstcount       => mm_interconnect_0_ram_uas_burstcount,    --      .burstcount
			uas_read             => mm_interconnect_0_ram_uas_read,          --      .read
			uas_write            => mm_interconnect_0_ram_uas_write,         --      .write
			uas_waitrequest      => mm_interconnect_0_ram_uas_waitrequest,   --      .waitrequest
			uas_readdatavalid    => mm_interconnect_0_ram_uas_readdatavalid, --      .readdatavalid
			uas_byteenable       => mm_interconnect_0_ram_uas_byteenable,    --      .byteenable
			uas_readdata         => mm_interconnect_0_ram_uas_readdata,      --      .readdata
			uas_writedata        => mm_interconnect_0_ram_uas_writedata,     --      .writedata
			uas_lock             => mm_interconnect_0_ram_uas_lock,          --      .lock
			uas_debugaccess      => mm_interconnect_0_ram_uas_debugaccess,   --      .debugaccess
			tcm_write_n_out      => ram_tcm_write_n_out,                     --   tcm.write_n_out
			tcm_read_out         => ram_tcm_read_out,                        --      .read_out
			tcm_chipselect_n_out => ram_tcm_chipselect_n_out,                --      .chipselect_n_out
			tcm_request          => ram_tcm_request,                         --      .request
			tcm_grant            => ram_tcm_grant,                           --      .grant
			tcm_address_out      => ram_tcm_address_out,                     --      .address_out
			tcm_data_out         => ram_tcm_data_out,                        --      .data_out
			tcm_data_outen       => ram_tcm_data_outen,                      --      .data_outen
			tcm_data_in          => ram_tcm_data_in                          --      .data_in
		);

	pin_sharer : component sopc_scope_sys_pin_sharer
		port map (
			clk_clk                  => clk_clk,                                     --   clk.clk
			reset_reset              => rst_controller_reset_out_reset,              -- reset.reset
			request                  => pin_sharer_tcm_request,                      --   tcm.request
			grant                    => pin_sharer_tcm_grant,                        --      .grant
			rom_tcm_read_out         => pin_sharer_tcm_rom_tcm_read_out_out,         --      .rom_tcm_read_out_out
			rom_tcm_chipselect_n_out => pin_sharer_tcm_rom_tcm_chipselect_n_out_out, --      .rom_tcm_chipselect_n_out_out
			ram_tcm_write_n_out      => pin_sharer_tcm_ram_tcm_write_n_out_out,      --      .ram_tcm_write_n_out_out
			ram_tcm_read_out         => pin_sharer_tcm_ram_tcm_read_out_out,         --      .ram_tcm_read_out_out
			ram_tcm_chipselect_n_out => pin_sharer_tcm_ram_tcm_chipselect_n_out_out, --      .ram_tcm_chipselect_n_out_out
			addr_out                 => pin_sharer_tcm_addr_out_out,                 --      .addr_out_out
			data_outen               => pin_sharer_tcm_data_outen_out,               --      .data_outen_out
			data_outen_in            => pin_sharer_tcm_data_outen_in,                --      .data_outen_in
			data_outen_outen         => pin_sharer_tcm_data_outen_outen,             --      .data_outen_outen
			tcs0_request             => ram_tcm_request,                             --  tcs0.request
			tcs0_grant               => ram_tcm_grant,                               --      .grant
			tcs0_address_out         => ram_tcm_address_out,                         --      .address_out
			tcs0_write_n_out(0)      => ram_tcm_write_n_out,                         --      .write_n_out
			tcs0_read_out(0)         => ram_tcm_read_out,                            --      .read_out
			tcs0_data_out            => ram_tcm_data_out,                            --      .data_out
			tcs0_data_in             => ram_tcm_data_in,                             --      .data_in
			tcs0_data_outen          => ram_tcm_data_outen,                          --      .data_outen
			tcs0_chipselect_n_out(0) => ram_tcm_chipselect_n_out,                    --      .chipselect_n_out
			tcs1_request             => rom_tcm_request,                             --  tcs1.request
			tcs1_grant               => rom_tcm_grant,                               --      .grant
			tcs1_address_out         => rom_tcm_address_out,                         --      .address_out
			tcs1_read_out(0)         => rom_tcm_read_out,                            --      .read_out
			tcs1_data_out            => rom_tcm_data_out,                            --      .data_out
			tcs1_data_in             => rom_tcm_data_in,                             --      .data_in
			tcs1_data_outen          => rom_tcm_data_outen,                          --      .data_outen
			tcs1_chipselect_n_out(0) => rom_tcm_chipselect_n_out                     --      .chipselect_n_out
		);

	bridge : component sopc_scope_sys_bridge
		port map (
			clk                          => clk_clk,                                     --   clk.clk
			reset                        => rst_controller_reset_out_reset,              -- reset.reset
			request                      => pin_sharer_tcm_request,                      --   tcs.request
			grant                        => pin_sharer_tcm_grant,                        --      .grant
			tcs_addr_out                 => pin_sharer_tcm_addr_out_out,                 --      .addr_out_out
			tcs_rom_tcm_chipselect_n_out => pin_sharer_tcm_rom_tcm_chipselect_n_out_out, --      .rom_tcm_chipselect_n_out_out
			tcs_ram_tcm_read_out         => pin_sharer_tcm_ram_tcm_read_out_out,         --      .ram_tcm_read_out_out
			tcs_ram_tcm_write_n_out      => pin_sharer_tcm_ram_tcm_write_n_out_out,      --      .ram_tcm_write_n_out_out
			tcs_data_outen               => pin_sharer_tcm_data_outen_out,               --      .data_outen_out
			tcs_data_outen_outen         => pin_sharer_tcm_data_outen_outen,             --      .data_outen_outen
			tcs_data_outen_in            => pin_sharer_tcm_data_outen_in,                --      .data_outen_in
			tcs_rom_tcm_read_out         => pin_sharer_tcm_rom_tcm_read_out_out,         --      .rom_tcm_read_out_out
			tcs_ram_tcm_chipselect_n_out => pin_sharer_tcm_ram_tcm_chipselect_n_out_out, --      .ram_tcm_chipselect_n_out_out
			addr_out                     => bridge_out_addr_out,                         --   out.addr_out
			rom_tcm_chipselect_n_out     => bridge_out_rom_tcm_chipselect_n_out,         --      .rom_tcm_chipselect_n_out
			ram_tcm_read_out             => bridge_out_ram_tcm_read_out,                 --      .ram_tcm_read_out
			ram_tcm_write_n_out          => bridge_out_ram_tcm_write_n_out,              --      .ram_tcm_write_n_out
			data_outen                   => bridge_out_data_outen,                       --      .data_outen
			rom_tcm_read_out             => bridge_out_rom_tcm_read_out,                 --      .rom_tcm_read_out
			ram_tcm_chipselect_n_out     => bridge_out_ram_tcm_chipselect_n_out          --      .ram_tcm_chipselect_n_out
		);

	rom : component sopc_scope_sys_rom
		generic map (
			TCM_ADDRESS_W                  => 19,
			TCM_DATA_W                     => 8,
			TCM_BYTEENABLE_W               => 1,
			TCM_READ_WAIT                  => 6,
			TCM_WRITE_WAIT                 => 0,
			TCM_SETUP_WAIT                 => 0,
			TCM_DATA_HOLD                  => 0,
			TCM_TURNAROUND_TIME            => 2,
			TCM_TIMING_UNITS               => 1,
			TCM_READLATENCY                => 2,
			TCM_SYMBOLS_PER_WORD           => 1,
			USE_READDATA                   => 1,
			USE_WRITEDATA                  => 1,
			USE_READ                       => 1,
			USE_WRITE                      => 0,
			USE_BYTEENABLE                 => 0,
			USE_CHIPSELECT                 => 1,
			USE_LOCK                       => 0,
			USE_ADDRESS                    => 1,
			USE_WAITREQUEST                => 0,
			USE_WRITEBYTEENABLE            => 0,
			USE_OUTPUTENABLE               => 0,
			USE_RESETREQUEST               => 0,
			USE_IRQ                        => 0,
			USE_RESET_OUTPUT               => 0,
			ACTIVE_LOW_READ                => 0,
			ACTIVE_LOW_LOCK                => 0,
			ACTIVE_LOW_WRITE               => 0,
			ACTIVE_LOW_CHIPSELECT          => 1,
			ACTIVE_LOW_BYTEENABLE          => 0,
			ACTIVE_LOW_OUTPUTENABLE        => 0,
			ACTIVE_LOW_WRITEBYTEENABLE     => 0,
			ACTIVE_LOW_WAITREQUEST         => 0,
			ACTIVE_LOW_BEGINTRANSFER       => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0
		)
		port map (
			clk_clk              => clk_clk,                                 --   clk.clk
			reset_reset          => rst_controller_reset_out_reset,          -- reset.reset
			uas_address          => mm_interconnect_0_rom_uas_address,       --   uas.address
			uas_burstcount       => mm_interconnect_0_rom_uas_burstcount,    --      .burstcount
			uas_read             => mm_interconnect_0_rom_uas_read,          --      .read
			uas_write            => mm_interconnect_0_rom_uas_write,         --      .write
			uas_waitrequest      => mm_interconnect_0_rom_uas_waitrequest,   --      .waitrequest
			uas_readdatavalid    => mm_interconnect_0_rom_uas_readdatavalid, --      .readdatavalid
			uas_byteenable       => mm_interconnect_0_rom_uas_byteenable,    --      .byteenable
			uas_readdata         => mm_interconnect_0_rom_uas_readdata,      --      .readdata
			uas_writedata        => mm_interconnect_0_rom_uas_writedata,     --      .writedata
			uas_lock             => mm_interconnect_0_rom_uas_lock,          --      .lock
			uas_debugaccess      => mm_interconnect_0_rom_uas_debugaccess,   --      .debugaccess
			tcm_read_out         => rom_tcm_read_out,                        --   tcm.read_out
			tcm_chipselect_n_out => rom_tcm_chipselect_n_out,                --      .chipselect_n_out
			tcm_request          => rom_tcm_request,                         --      .request
			tcm_grant            => rom_tcm_grant,                           --      .grant
			tcm_address_out      => rom_tcm_address_out,                     --      .address_out
			tcm_data_out         => rom_tcm_data_out,                        --      .data_out
			tcm_data_outen       => rom_tcm_data_outen,                      --      .data_outen
			tcm_data_in          => rom_tcm_data_in                          --      .data_in
		);

	mm_interconnect_0 : component sopc_scope_sys_mm_interconnect_0
		port map (
			clk_0_clk_clk                            => clk_clk,                                              --                          clk_0_clk.clk
			nios_reset_n_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                       -- nios_reset_n_reset_bridge_in_reset.reset
			nios_data_master_address                 => nios_data_master_address,                             --                   nios_data_master.address
			nios_data_master_waitrequest             => nios_data_master_waitrequest,                         --                                   .waitrequest
			nios_data_master_byteenable              => nios_data_master_byteenable,                          --                                   .byteenable
			nios_data_master_read                    => nios_data_master_read,                                --                                   .read
			nios_data_master_readdata                => nios_data_master_readdata,                            --                                   .readdata
			nios_data_master_readdatavalid           => nios_data_master_readdatavalid,                       --                                   .readdatavalid
			nios_data_master_write                   => nios_data_master_write,                               --                                   .write
			nios_data_master_writedata               => nios_data_master_writedata,                           --                                   .writedata
			nios_data_master_debugaccess             => nios_data_master_debugaccess,                         --                                   .debugaccess
			nios_instruction_master_address          => nios_instruction_master_address,                      --            nios_instruction_master.address
			nios_instruction_master_waitrequest      => nios_instruction_master_waitrequest,                  --                                   .waitrequest
			nios_instruction_master_read             => nios_instruction_master_read,                         --                                   .read
			nios_instruction_master_readdata         => nios_instruction_master_readdata,                     --                                   .readdata
			nios_instruction_master_readdatavalid    => nios_instruction_master_readdatavalid,                --                                   .readdatavalid
			jtag_avalon_jtag_slave_address           => mm_interconnect_0_jtag_avalon_jtag_slave_address,     --             jtag_avalon_jtag_slave.address
			jtag_avalon_jtag_slave_write             => mm_interconnect_0_jtag_avalon_jtag_slave_write,       --                                   .write
			jtag_avalon_jtag_slave_read              => mm_interconnect_0_jtag_avalon_jtag_slave_read,        --                                   .read
			jtag_avalon_jtag_slave_readdata          => mm_interconnect_0_jtag_avalon_jtag_slave_readdata,    --                                   .readdata
			jtag_avalon_jtag_slave_writedata         => mm_interconnect_0_jtag_avalon_jtag_slave_writedata,   --                                   .writedata
			jtag_avalon_jtag_slave_waitrequest       => mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest, --                                   .waitrequest
			jtag_avalon_jtag_slave_chipselect        => mm_interconnect_0_jtag_avalon_jtag_slave_chipselect,  --                                   .chipselect
			nios_jtag_debug_module_address           => mm_interconnect_0_nios_jtag_debug_module_address,     --             nios_jtag_debug_module.address
			nios_jtag_debug_module_write             => mm_interconnect_0_nios_jtag_debug_module_write,       --                                   .write
			nios_jtag_debug_module_read              => mm_interconnect_0_nios_jtag_debug_module_read,        --                                   .read
			nios_jtag_debug_module_readdata          => mm_interconnect_0_nios_jtag_debug_module_readdata,    --                                   .readdata
			nios_jtag_debug_module_writedata         => mm_interconnect_0_nios_jtag_debug_module_writedata,   --                                   .writedata
			nios_jtag_debug_module_byteenable        => mm_interconnect_0_nios_jtag_debug_module_byteenable,  --                                   .byteenable
			nios_jtag_debug_module_waitrequest       => mm_interconnect_0_nios_jtag_debug_module_waitrequest, --                                   .waitrequest
			nios_jtag_debug_module_debugaccess       => mm_interconnect_0_nios_jtag_debug_module_debugaccess, --                                   .debugaccess
			ram_uas_address                          => mm_interconnect_0_ram_uas_address,                    --                            ram_uas.address
			ram_uas_write                            => mm_interconnect_0_ram_uas_write,                      --                                   .write
			ram_uas_read                             => mm_interconnect_0_ram_uas_read,                       --                                   .read
			ram_uas_readdata                         => mm_interconnect_0_ram_uas_readdata,                   --                                   .readdata
			ram_uas_writedata                        => mm_interconnect_0_ram_uas_writedata,                  --                                   .writedata
			ram_uas_burstcount                       => mm_interconnect_0_ram_uas_burstcount,                 --                                   .burstcount
			ram_uas_byteenable                       => mm_interconnect_0_ram_uas_byteenable,                 --                                   .byteenable
			ram_uas_readdatavalid                    => mm_interconnect_0_ram_uas_readdatavalid,              --                                   .readdatavalid
			ram_uas_waitrequest                      => mm_interconnect_0_ram_uas_waitrequest,                --                                   .waitrequest
			ram_uas_lock                             => mm_interconnect_0_ram_uas_lock,                       --                                   .lock
			ram_uas_debugaccess                      => mm_interconnect_0_ram_uas_debugaccess,                --                                   .debugaccess
			rom_uas_address                          => mm_interconnect_0_rom_uas_address,                    --                            rom_uas.address
			rom_uas_write                            => mm_interconnect_0_rom_uas_write,                      --                                   .write
			rom_uas_read                             => mm_interconnect_0_rom_uas_read,                       --                                   .read
			rom_uas_readdata                         => mm_interconnect_0_rom_uas_readdata,                   --                                   .readdata
			rom_uas_writedata                        => mm_interconnect_0_rom_uas_writedata,                  --                                   .writedata
			rom_uas_burstcount                       => mm_interconnect_0_rom_uas_burstcount,                 --                                   .burstcount
			rom_uas_byteenable                       => mm_interconnect_0_rom_uas_byteenable,                 --                                   .byteenable
			rom_uas_readdatavalid                    => mm_interconnect_0_rom_uas_readdatavalid,              --                                   .readdatavalid
			rom_uas_waitrequest                      => mm_interconnect_0_rom_uas_waitrequest,                --                                   .waitrequest
			rom_uas_lock                             => mm_interconnect_0_rom_uas_lock,                       --                                   .lock
			rom_uas_debugaccess                      => mm_interconnect_0_rom_uas_debugaccess,                --                                   .debugaccess
			temp_ram_s1_address                      => mm_interconnect_0_temp_ram_s1_address,                --                        temp_ram_s1.address
			temp_ram_s1_write                        => mm_interconnect_0_temp_ram_s1_write,                  --                                   .write
			temp_ram_s1_readdata                     => mm_interconnect_0_temp_ram_s1_readdata,               --                                   .readdata
			temp_ram_s1_writedata                    => mm_interconnect_0_temp_ram_s1_writedata,              --                                   .writedata
			temp_ram_s1_chipselect                   => mm_interconnect_0_temp_ram_s1_chipselect,             --                                   .chipselect
			temp_ram_s1_clken                        => mm_interconnect_0_temp_ram_s1_clken                   --                                   .clken
		);

	irq_mapper : component sopc_scope_sys_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			sender_irq    => nios_d_irq_irq                  --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios_jtag_debug_module_reset_reset, -- reset_in0.reset
			reset_in1      => nios_jtag_debug_module_reset_reset, -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_avalon_jtag_slave_write;

	mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_avalon_jtag_slave_read;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of sopc_scope_sys
